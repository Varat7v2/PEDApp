*Generated netlist for the circuit diagram.
L1 2 3 120
V1 1 0 21
C1 3 0 577
D1 2 0 1N4148
R2 4 0 0.8485547322214142
.lib /home/varat/Documents/LTspiceXVII/lib/cmp/standard.dio
.options TEMP = 25C
.options TNOM = 25C
.tran 100m
.model switch SW(Ron=1m Roff=100Meg Vt=0.5 Vh=0)
.end