*Generated netlist for the circuit diagram.
L1 0 0 104
V1 0 0 45
C1 0 0 627
D1 0 0 1N4148
R2 0 0 1.06
.libraries /home/varat/Documents/LTspiceXVII/libraries/cmp/standard.dio
.options TEMP = 25C
.options TNOM = 25C
.tran 100m
.model switch SW(Ron=1m Roff=100Meg Vt=0.5 Vh=0)
.end